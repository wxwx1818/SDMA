`ifndef _NSDM_VH
`define _NSDM_VH

// +[1] DEFINE Design Version DECLARATION (XJB)----------------------------------------------------------------------------------------------------
`define		HIGH_BANDWIDTH_VERSION
// `define		MED_BADNWIDTH_VERSION
// +[1] DEFINE Design Version DECLARATION----------------------------------------------------------------------------------------------------

// +[2] DEFINE NSDM GMV Inout Port DECLARATION (WX)----------------------------------------------------------------------------------------------------
// ++About address width--------------------------------------------------
`define		SDMA_ADDRWIDTH								32
// ++About cache data width--------------------------------------------------
`define		SDMA_CACHEDATAWIDTH							512
// ++About ahb data width--------------------------------------------------
`ifdef HIGH_BANDWIDTH_VERSION		
	`define	SDMA_AHBDATAWIDTH							128
`else		
`ifdef MED_BADNWIDTH_VERSION 		
	`define	SDMA_AHBDATAWIDTH							64
`else		
	`define SDMA_AHBDATAWIDTH							32	
`endif		
`endif		
`define SDMA_SECTION_DINNUMDATAWIDTH					$clog2(`SDMA_CACHEDATAWIDTH/8)+1		//bytes number
// -[2] DEFINE NSDM GMV Inout Port DECLARATION----------------------------------------------------------------------------------------------------

// +[3] DEFINE NMD Macro Instruction DECLARATION (WX)----------------------------------------------------------------------------------------------------
`define	SDMA_INSTWIDTH						640

`define SDMA_INST_SDMAMODESTART				0
`define SDMA_INST_SDMAMODEWIDTH				6
`define SDMA_INST_SDMAMODEEND				`SDMA_INST_SDMAMODESTART + `SDMA_INST_SDMAMODEWIDTH - 1

`define SDMA_INST_SRCPORTIDSTART			`SDMA_INST_SDMAMODEEND + 1
`define SDMA_INST_SRCPORTIDWIDTH			3
`define SDMA_INST_SRCPORTIDEND				`SDMA_INST_SRCPORTIDSTART + `SDMA_INST_SRCPORTIDWIDTH - 1

`define SDMA_INST_DSTPORTIDSTART			`SDMA_INST_SRCPORTIDEND + 1
`define SDMA_INST_DSTPORTIDWIDTH			3
`define SDMA_INST_DSTPORTIDEND				`SDMA_INST_DSTPORTIDSTART + `SDMA_INST_DSTPORTIDWIDTH - 1

`define SDMA_INST_SRCFMSADDRSTART			`SDMA_INST_DSTPORTIDEND + 1
`define SDMA_INST_SRCFMSADDRWIDTH			32
`define SDMA_INST_SRCFMSADDREND				`SDMA_INST_SRCFMSADDRSTART + `SDMA_INST_SRCFMSADDRWIDTH - 1

`define SDMA_INST_DSTFMSADDRSTART			`SDMA_INST_SRCFMSADDREND + 1
`define SDMA_INST_DSTFMSADDRWIDTH			32
`define SDMA_INST_DSTFMSADDREND				`SDMA_INST_DSTFMSADDRSTART + `SDMA_INST_DSTFMSADDRWIDTH - 1

`define SDMA_INST_SRCFMSMOVELENGTHSTART		`SDMA_INST_DSTFMSADDREND + 1
`define SDMA_INST_SRCFMSMOVELENGTHWIDTH		21
`define SDMA_INST_SRCFMSMOVELENGTHEND		`SDMA_INST_SRCFMSMOVELENGTHSTART + `SDMA_INST_SRCFMSMOVELENGTHWIDTH - 1

`define SDMA_INST_SRCFMS2ADDRSTART			`SDMA_INST_SRCFMSMOVELENGTHEND + 1
`define SDMA_INST_SRCFMS2ADDRWIDTH			32
`define SDMA_INST_SRCFMS2ADDREND			`SDMA_INST_SRCFMS2ADDRSTART + `SDMA_INST_SRCFMS2ADDRWIDTH - 1

`define SDMA_INST_SRCFMS1CONCATELENGTHSTART	`SDMA_INST_SRCFMS2ADDREND + 1
`define SDMA_INST_SRCFMS1CONCATELENGTHWIDTH	21
`define SDMA_INST_SRCFMS1CONCATELENGTHEND	`SDMA_INST_SRCFMS1CONCATELENGTHSTART + `SDMA_INST_SRCFMS1CONCATELENGTHWIDTH - 1

`define SDMA_INST_SRCFMS2CONCATELENGTHSTART	`SDMA_INST_SRCFMS1CONCATELENGTHEND + 1
`define SDMA_INST_SRCFMS2CONCATELENGTHWIDTH	21
`define SDMA_INST_SRCFMS2CONCATELENGTHEND	`SDMA_INST_SRCFMS2CONCATELENGTHSTART + `SDMA_INST_SRCFMS2CONCATELENGTHWIDTH - 1

`define SDMA_INST_SRCFMS2MOVELENGTHSTART	`SDMA_INST_SRCFMS2CONCATELENGTHEND + 1
`define SDMA_INST_SRCFMS2MOVELENGTHWIDTH	21
`define SDMA_INST_SRCFMS2MOVELENGTHEND		`SDMA_INST_SRCFMS2MOVELENGTHSTART + `SDMA_INST_SRCFMS2MOVELENGTHWIDTH - 1

`define SDMA_INST_SRCFMSCSTART				`SDMA_INST_SRCFMS2MOVELENGTHEND + 1
`define SDMA_INST_SRCFMSCWIDTH				13
`define SDMA_INST_SRCFMSCEND				`SDMA_INST_SRCFMSCSTART + `SDMA_INST_SRCFMSCWIDTH - 1

`define SDMA_INST_SRCFMSXSTART				`SDMA_INST_SRCFMSCEND + 1
`define SDMA_INST_SRCFMSXWIDTH				13
`define SDMA_INST_SRCFMSXEND				`SDMA_INST_SRCFMSXSTART + `SDMA_INST_SRCFMSXWIDTH - 1

`define SDMA_INST_SRCFMSYSTART				`SDMA_INST_SRCFMSXEND + 1
`define SDMA_INST_SRCFMSYWIDTH				13
`define SDMA_INST_SRCFMSYEND				`SDMA_INST_SRCFMSYSTART + `SDMA_INST_SRCFMSYWIDTH - 1

`define SDMA_INST_DSTFMSSTRIDE3START		`SDMA_INST_SRCFMSYEND + 1
`define SDMA_INST_DSTFMSSTRIDE3WIDTH		17
`define SDMA_INST_DSTFMSSTRIDE3END			`SDMA_INST_DSTFMSSTRIDE3START + `SDMA_INST_DSTFMSSTRIDE3WIDTH - 1

`define SDMA_INST_DSTFMSSTRIDE2START		`SDMA_INST_DSTFMSSTRIDE3END + 1
`define SDMA_INST_DSTFMSSTRIDE2WIDTH		17
`define SDMA_INST_DSTFMSSTRIDE2END			`SDMA_INST_DSTFMSSTRIDE2START + `SDMA_INST_DSTFMSSTRIDE2WIDTH - 1

`define SDMA_INST_DSTFMSSTRIDE1START		`SDMA_INST_DSTFMSSTRIDE2END + 1
`define SDMA_INST_DSTFMSSTRIDE1WIDTH		17
`define SDMA_INST_DSTFMSSTRIDE1END			`SDMA_INST_DSTFMSSTRIDE1START + `SDMA_INST_DSTFMSSTRIDE1WIDTH - 1

`define SDMA_INST_PADDINGAXISBEFORESTART	`SDMA_INST_DSTFMSSTRIDE1END + 1
`define SDMA_INST_PADDINGAXISBEFOREWIDTH	3
`define SDMA_INST_PADDINGAXISBEFOREEND		`SDMA_INST_PADDINGAXISBEFORESTART + `SDMA_INST_PADDINGAXISBEFOREWIDTH - 1

`define SDMA_INST_PADDINGLEFTXSTART			`SDMA_INST_PADDINGAXISBEFOREEND + 1
`define SDMA_INST_PADDINGLEFTXWIDTH			6
`define SDMA_INST_PADDINGLEFTXEND			`SDMA_INST_PADDINGLEFTXSTART + `SDMA_INST_PADDINGLEFTXWIDTH - 1

`define SDMA_INST_PADDINGRIGHTXSTART		`SDMA_INST_PADDINGLEFTXEND + 1
`define SDMA_INST_PADDINGRIGHTXWIDTH		6
`define SDMA_INST_PADDINGRIGHTXEND			`SDMA_INST_PADDINGRIGHTXSTART + `SDMA_INST_PADDINGRIGHTXWIDTH - 1

`define SDMA_INST_PADDINGLEFTYSTART			`SDMA_INST_PADDINGRIGHTXEND + 1
`define SDMA_INST_PADDINGLEFTYWIDTH			6
`define SDMA_INST_PADDINGLEFTYEND			`SDMA_INST_PADDINGLEFTYSTART + `SDMA_INST_PADDINGLEFTYWIDTH - 1

`define SDMA_INST_PADDINGRIGHTYSTART		`SDMA_INST_PADDINGLEFTYEND + 1
`define SDMA_INST_PADDINGRIGHTYWIDTH		6
`define SDMA_INST_PADDINGRIGHTYEND			`SDMA_INST_PADDINGRIGHTYSTART + `SDMA_INST_PADDINGRIGHTYWIDTH - 1

`define SDMA_INST_INSERTZERONUMSTART		`SDMA_INST_PADDINGRIGHTYEND + 1
`define SDMA_INST_INSERTZERONUMWIDTH		3
`define SDMA_INST_INSERTZERONUMEND			`SDMA_INST_INSERTZERONUMSTART + `SDMA_INST_INSERTZERONUMWIDTH - 1

`define SDMA_INST_INSERTZERONUMTOTALXSTART	`SDMA_INST_INSERTZERONUMEND + 1
`define SDMA_INST_INSERTZERONUMTOTALXWIDTH	11
`define SDMA_INST_INSERTZERONUMTOTALXEND	`SDMA_INST_INSERTZERONUMTOTALXSTART + `SDMA_INST_INSERTZERONUMTOTALXWIDTH - 1

`define SDMA_INST_INSERTZERONUMTOTALYSTART	`SDMA_INST_INSERTZERONUMTOTALXEND + 1
`define SDMA_INST_INSERTZERONUMTOTALYWIDTH	11
`define SDMA_INST_INSERTZERONUMTOTALYEND	`SDMA_INST_INSERTZERONUMTOTALYSTART + `SDMA_INST_INSERTZERONUMTOTALYWIDTH - 1

`define SDMA_INST_UPSAMPLEIDXXSTART			`SDMA_INST_INSERTZERONUMTOTALYEND + 1
`define SDMA_INST_UPSAMPLEIDXXWIDTH			3
`define SDMA_INST_UPSAMPLEIDXXEND			`SDMA_INST_UPSAMPLEIDXXSTART + `SDMA_INST_UPSAMPLEIDXXWIDTH - 1

`define SDMA_INST_UPSAMPLEIDXYSTART			`SDMA_INST_UPSAMPLEIDXXEND + 1
`define SDMA_INST_UPSAMPLEIDXYWIDTH			3
`define SDMA_INST_UPSAMPLEIDXYEND			`SDMA_INST_UPSAMPLEIDXYSTART + `SDMA_INST_UPSAMPLEIDXYWIDTH - 1

`define SDMA_INST_CROPFMSSTRIDE2START		`SDMA_INST_UPSAMPLEIDXYEND + 1
`define SDMA_INST_CROPFMSSTRIDE2WIDTH		17
`define SDMA_INST_CROPFMSSTRIDE2END			`SDMA_INST_CROPFMSSTRIDE2START + `SDMA_INST_CROPFMSSTRIDE2WIDTH - 1

`define SDMA_INST_CROPFMSSTRIDE1START		`SDMA_INST_CROPFMSSTRIDE2END + 1
`define SDMA_INST_CROPFMSSTRIDE1WIDTH		13
`define SDMA_INST_CROPFMSSTRIDE1END			`SDMA_INST_CROPFMSSTRIDE1START + `SDMA_INST_CROPFMSSTRIDE1WIDTH - 1

`define SDMA_INST_CROPFMSCSTART				`SDMA_INST_CROPFMSSTRIDE1END + 1
`define SDMA_INST_CROPFMSCWIDTH				13
`define SDMA_INST_CROPFMSCEND				`SDMA_INST_CROPFMSCSTART + `SDMA_INST_CROPFMSCWIDTH - 1

`define SDMA_INST_CROPFMSXSTART				`SDMA_INST_CROPFMSCEND + 1
`define SDMA_INST_CROPFMSXWIDTH				13
`define SDMA_INST_CROPFMSXEND				`SDMA_INST_CROPFMSXSTART + `SDMA_INST_CROPFMSXWIDTH - 1

`define SDMA_INST_CROPFMSYSTART				`SDMA_INST_CROPFMSXEND + 1
`define SDMA_INST_CROPFMSYWIDTH				13
`define SDMA_INST_CROPFMSYEND				`SDMA_INST_CROPFMSYSTART + `SDMA_INST_CROPFMSYWIDTH - 1

`define SDMA_INST_CROPFMS2STRIDE2START		`SDMA_INST_CROPFMSYEND + 1
`define SDMA_INST_CROPFMS2STRIDE2WIDTH		17
`define SDMA_INST_CROPFMS2STRIDE2END		`SDMA_INST_CROPFMS2STRIDE2START + `SDMA_INST_CROPFMS2STRIDE2WIDTH - 1

`define SDMA_INST_CROPFMS2STRIDE1START		`SDMA_INST_CROPFMS2STRIDE2END + 1
`define SDMA_INST_CROPFMS2STRIDE1WIDTH		13
`define SDMA_INST_CROPFMS2STRIDE1END		`SDMA_INST_CROPFMS2STRIDE1START + `SDMA_INST_CROPFMS2STRIDE1WIDTH - 1

`define SDMA_INST_CROPFMS2CSTART			`SDMA_INST_CROPFMS2STRIDE1END + 1
`define SDMA_INST_CROPFMS2CWIDTH			13
`define SDMA_INST_CROPFMS2CEND				`SDMA_INST_CROPFMS2CSTART + `SDMA_INST_CROPFMS2CWIDTH - 1

`define SDMA_INST_CROPFMS2XSTART			`SDMA_INST_CROPFMS2CEND + 1
`define SDMA_INST_CROPFMS2XWIDTH			13
`define SDMA_INST_CROPFMS2XEND				`SDMA_INST_CROPFMS2XSTART + `SDMA_INST_CROPFMS2XWIDTH - 1

`define SDMA_INST_CROPFMS2YSTART			`SDMA_INST_CROPFMS2XEND + 1
`define SDMA_INST_CROPFMS2YWIDTH			13
`define SDMA_INST_CROPFMS2YEND				`SDMA_INST_CROPFMS2YSTART + `SDMA_INST_CROPFMS2YWIDTH - 1

`define SDMA_INST_SRCFMSCYCSADDRSTART		`SDMA_INST_CROPFMS2YEND + 1
`define SDMA_INST_SRCFMSCYCSADDRWIDTH		32
`define SDMA_INST_SRCFMSCYCSADDREND			`SDMA_INST_SRCFMSCYCSADDRSTART + `SDMA_INST_SRCFMSCYCSADDRWIDTH - 1

`define SDMA_INST_SRCFMSCYCEADDRSTART		`SDMA_INST_SRCFMSCYCSADDREND + 1
`define	SDMA_INST_SRCFMSCYCEADDRWIDTH		32
`define SDMA_INST_SRCFMSCYCEADDREND			`SDMA_INST_SRCFMSCYCEADDRSTART + `SDMA_INST_SRCFMSCYCEADDRWIDTH - 1

`define SDMA_INST_SRCFMSCYCALIGNENASTART	`SDMA_INST_SRCFMSCYCEADDREND + 1
`define SDMA_INST_SRCFMSCYCALIGNENAWIDTH	1
`define SDMA_INST_SRCFMSCYCALIGNENAEND		`SDMA_INST_SRCFMSCYCALIGNENASTART + `SDMA_INST_SRCFMSCYCALIGNENAWIDTH - 1
// -[3] DEFINE NSDM GMV Macro Instruction DECLARATION----------------------------------------------------------------------------------------------------

// +[4] DEFINE NSDM GMV Transfer Mode DECLARATION (WX)----------------------------------------------------------------------------------------------------
// Try to avoid AHB nonseq write as much as possiable.

`define	SDMA_SDP_MODE_AHB2AHBSEQ		   		0			//src: 32b  valid/write  dst: 32b  valid/read
`define	SDMA_SDP_MODE_AHB2AHBNONSEQ     		1			//src: 32b  valid/write	 dst: 8b   valid/read
`define SDMA_SDP_MODE_AHB2CACHESEQ				2			//src: 32b  valid/write  dst: 512b valid/read
`define	SDMA_SDP_MODE_AHB2CACHENONSEQ   		3			//src: 32b  valid/write  dst: 8b   valid/read
`define SDMA_SDP_MODE_CACHE2AHBSEQ 	   			4			//src: 512b valid/write	 dst: 32b  valid/read
`define SDMA_SDP_MODE_CACHE2AHBNONSEQ   		5			//src: 512b valid/write	 dst: 8b   valid/read
`define SDMA_SDP_MODE_CACHE2CACHESEQ	   		6			//src: 512b valid/write  dst: 512b valid/read
`define SDMA_SDP_MODE_CACHE2CACHENONSEQ 		7			//src: 512b valid/write	 dst: 8b   valid/read
// -[4] DEFINE NSDM GMV Transfer Mode DECLARATION----------------------------------------------------------------------------------------------------

// +[5] DEFINE NSDM NMV Width DECLARATION (XJB)----------------------------------------------------------------------------------------------------
`define 	NMV_PARAM_ADDR_WIDTH						32
`define 	NMV_PARAM_NUM_WIDTH							16
`define 	NMV_INSTR_ADDR_WIDTH						`NMV_PARAM_ADDR_WIDTH
`define 	NMV_INSTR_NUM_WIDTH							`NMV_PARAM_NUM_WIDTH
// -[5] DEFINE NSDM NMV Width DECLARATION----------------------------------------------------------------------------------------------------

`endif // _NSDM_VH
